/******************************************************************************
* SPECT - DPI
*
* TODO: License
*
* Author: Marek Santa
******************************************************************************/
`ifndef SPECT_ISS_DPI_TYPES_SVH
`define SPECT_ISS_DPI_TYPES_SVH


/////////////////////////////////////////////////////////////////////////////
// Typedefs
/////////////////////////////////////////////////////////////////////////////
typedef enum {
  DPI_SPECT_DATA_RAM_IN       = (1 << 0),
  DPI_SPECT_DATA_RAM_OUT      = (1 << 1),
  DPI_SPECT_CONST_ROM         = (1 << 2),
  DPI_SPECT_INSTRUCTION_MEM   = (1 << 3)
} dpi_mem_type_t;

typedef enum {
  DPI_SPECT_FLAG_ZERO         = (1 << 0),
  DPI_SPECT_FLAG_CARRY        = (1 << 1)
} dpi_flag_type_t;

typedef enum {
  DPI_SPECT_INT_DONE          = (1 << 0),
  DPI_SPECT_INT_ERR           = (1 << 1)
} dpi_int_type_t;

typedef enum {
  DPI_CHANGE_GPR              = (1 << 0),
  DPI_CHANGE_FLAG             = (1 << 1),
  DPI_CHANGE_MEM              = (1 << 2),
  DPI_CHANGE_SRR              = (1 << 3),
  DPI_CHANGE_INT              = (1 << 4),
  DPI_CHANGE_RAR              = (1 << 5),
  DPI_CHANGE_RAR_SP           = (1 << 6)
} dpi_change_kind_t;

typedef struct {
    dpi_change_kind_t kind;

    // Identifies object on which change occured based on kind
    //  DPI_CHANGE_GPR:
    //      0  - GPR0
    //      ...
    //      31 - GPR31
    //
    //  DPI_CHANGE_FLAG:
    //      DPI_SPECT_FLAG_ZERO
    //      DPI_SPECT_FLAG_CARRY
    //
    //  DPI_CHANGE_MEM:
    //      Address in memory on which change occured.
    //
    //  DPI_CHANGE_SRR:
    //      -
    //
    //  DPI_CHANGE_INT:
    //      DPI_SPECT_INT_DONE
    //      DPI_SPECT_INT_ERR
    //
    //  DPI_CHANGE_RAR:
    //      0 - G_RAR_DEPTH - Index of RAR stack where changed occured
    //
    //  DPI_CAHNGE_RAR_SP:
    //      -
    int               obj;

    // Old / New value of the object based  on 'kind':
    //  DPI_CHANGE_GPR:
    //      0 - Bits 31:0
    //      ...
    //      7 - Bits 255:232
    //
    //  DPI_CHANGE_FLAG:
    //      0 - Value of flag
    //
    //  DPI_CHANGE_MEM:
    //      0 - Bits 31:0 of memory location
    //
    //  DPI_CHANGE_INT:
    //      0 - Value of the interrupt
    //
    //  DPI_CHANGE_RAR:
    //      0 - Bits 31:0 of RAR stack location
    //
    //  DPI_CAHNGE_RAR_SP:
    //      Value of RAR stack pointer
    int               old_val[8];
    int               new_val[8];
} dpi_state_change_t;

`endif // SPECT_ISS_DPI_TYPES_SVH
